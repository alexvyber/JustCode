module main

fn main() {
    i := 0
    x := 1

    println(x)
    }
