

module module_long_name_here_goes

pub fn hi() {
    println('hi form long')
    }
