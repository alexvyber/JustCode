module main

fn main () {

    a := false 

    if a {
        println("true")
        } else {
            println("false")
            }



        }
