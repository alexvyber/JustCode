module main

const b = 3
fn main () {
println(b)
println(a)
println(take)
}

fn return3 () int { return 3 }

const take = return3()


const a = 4

